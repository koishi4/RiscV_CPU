`include "defines.vh"

module ex_stage(
    input clk,
    input rst_n
);
    // TODO: execute/ALU stage.
endmodule
