`include "defines.vh"

module trap_ctrl(
    input clk,
    input rst_n
);
    // TODO: trap entry/return control (mret).
endmodule
