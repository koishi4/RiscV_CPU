module mem_model;
    // TODO: optional behavioral memory model for testbench.
endmodule
