`timescale 1ns/1ps
`include "defines.vh"
`include "interface.vh"

module cpu_top(
    input  clk,
    input  rst_n,
    `MEM_REQ_PORTS(output, cpu_mem),
    `MEM_RSP_PORTS(input, cpu_mem),
    `MULDIV_REQ_PORTS(output, muldiv),
    `MULDIV_RSP_PORTS(input, muldiv),
    input  ext_irq
);
    // TODO: implement 2-hart RV32 core, CSR/trap, and muldiv integration.
    reg [`HART_NUM-1:0] blocked;
    reg [`HART_NUM-1:0] blocked_n;
    reg [`XLEN-1:0] pc[`HART_NUM-1:0];
    reg ifid_valid[`HART_NUM-1:0];
    reg [`XLEN-1:0] ifid_pc[`HART_NUM-1:0];
    reg [31:0] ifid_inst[`HART_NUM-1:0];
    reg idex_valid[`HART_NUM-1:0];
    reg [`XLEN-1:0] idex_pc[`HART_NUM-1:0];
    reg [31:0] idex_inst[`HART_NUM-1:0];
    reg [`HART_ID_W-1:0] idex_hart_id[`HART_NUM-1:0];
    reg [`REG_ADDR_W-1:0] idex_rs1[`HART_NUM-1:0];
    reg [`REG_ADDR_W-1:0] idex_rs2[`HART_NUM-1:0];
    reg [`REG_ADDR_W-1:0] idex_rd[`HART_NUM-1:0];
    reg [6:0] idex_opcode[`HART_NUM-1:0];
    reg [2:0] idex_funct3[`HART_NUM-1:0];
    reg [6:0] idex_funct7[`HART_NUM-1:0];
    reg [`XLEN-1:0] idex_imm[`HART_NUM-1:0];
    reg [`XLEN-1:0] idex_rs1_val[`HART_NUM-1:0];
    reg [`XLEN-1:0] idex_rs2_val[`HART_NUM-1:0];
    reg exmem_valid[`HART_NUM-1:0];
    reg [`HART_ID_W-1:0] exmem_hart_id[`HART_NUM-1:0];
    reg [`REG_ADDR_W-1:0] exmem_rd[`HART_NUM-1:0];
    reg [`XLEN-1:0] exmem_alu_result[`HART_NUM-1:0];
    reg [`XLEN-1:0] exmem_rs2_val[`HART_NUM-1:0];
    reg exmem_is_load[`HART_NUM-1:0];
    reg exmem_mem_we[`HART_NUM-1:0];
    reg exmem_wb_en[`HART_NUM-1:0];
    reg [`XLEN-1:0] exmem_wb_data_raw[`HART_NUM-1:0];
    reg exwb_valid[`HART_NUM-1:0];
    reg [`HART_ID_W-1:0] exwb_hart_id[`HART_NUM-1:0];
    reg [`REG_ADDR_W-1:0] exwb_rd[`HART_NUM-1:0];
    reg [`XLEN-1:0] exwb_data[`HART_NUM-1:0];
    reg muldiv_pending;
    reg [`XLEN-1:0] muldiv_pending_result;
    reg [`HART_ID_W-1:0] muldiv_pending_hart_id;
    reg [`REG_ADDR_W-1:0] muldiv_pending_rd;
    reg [`HART_ID_W-1:0] ifetch_hart_d;
    reg [`XLEN-1:0] ifetch_pc_d;
    reg ifetch_req;
    reg mem_inflight;
    reg mem_inflight_is_data;
    reg [`ADDR_W-1:0] mem_inflight_addr;
    reg mem_inflight_we;
    reg [`XLEN-1:0] mem_inflight_wdata;
    reg ifetch_kill[`HART_NUM-1:0];
    reg mem_req_d;
    reg mem_is_data_d;
    integer h;

    wire [`HART_ID_W-1:0] cur_hart;
    wire cur_valid;
    wire [`HART_ID_W-1:0] exec_hart = cur_hart;
    wire exec_valid = cur_valid;

    wire ifid_valid_cur = ifid_valid[exec_hart];
    wire [`XLEN-1:0] ifid_pc_cur = ifid_pc[exec_hart];
    wire [31:0] ifid_inst_cur = ifid_inst[exec_hart];
    wire idex_valid_cur = idex_valid[exec_hart];
    wire [`XLEN-1:0] idex_pc_cur = idex_pc[exec_hart];
    wire [31:0] idex_inst_cur = idex_inst[exec_hart];
    wire [`HART_ID_W-1:0] idex_hart_id_cur = idex_hart_id[exec_hart];
    wire [`REG_ADDR_W-1:0] idex_rs1_cur = idex_rs1[exec_hart];
    wire [`REG_ADDR_W-1:0] idex_rs2_cur = idex_rs2[exec_hart];
    wire [`REG_ADDR_W-1:0] idex_rd_cur = idex_rd[exec_hart];
    wire [6:0] idex_opcode_cur = idex_opcode[exec_hart];
    wire [2:0] idex_funct3_cur = idex_funct3[exec_hart];
    wire [6:0] idex_funct7_cur = idex_funct7[exec_hart];
    wire [`XLEN-1:0] idex_imm_cur = idex_imm[exec_hart];
    wire [`XLEN-1:0] idex_rs1_val_cur = idex_rs1_val[exec_hart];
    wire [`XLEN-1:0] idex_rs2_val_cur = idex_rs2_val[exec_hart];
    wire exmem_valid_cur = exmem_valid[exec_hart];
    wire [`HART_ID_W-1:0] exmem_hart_id_cur = exmem_hart_id[exec_hart];
    wire [`REG_ADDR_W-1:0] exmem_rd_cur = exmem_rd[exec_hart];
    wire [`XLEN-1:0] exmem_alu_result_cur = exmem_alu_result[exec_hart];
    wire [`XLEN-1:0] exmem_rs2_val_cur = exmem_rs2_val[exec_hart];
    wire exmem_is_load_cur = exmem_is_load[exec_hart];
    wire exmem_mem_we_cur = exmem_mem_we[exec_hart];
    wire exmem_wb_en_cur = exmem_wb_en[exec_hart];
    wire [`XLEN-1:0] exmem_wb_data_raw_cur = exmem_wb_data_raw[exec_hart];
    wire exwb_valid_cur = exwb_valid[exec_hart];
    wire [`HART_ID_W-1:0] exwb_hart_id_cur = exwb_hart_id[exec_hart];
    wire [`REG_ADDR_W-1:0] exwb_rd_cur = exwb_rd[exec_hart];
    wire [`XLEN-1:0] exwb_data_cur = exwb_data[exec_hart];

    wire [`REG_ADDR_W-1:0] raddr1 = ifid_valid_cur ? ifid_inst_cur[19:15] : {`REG_ADDR_W{1'b0}};
    wire [`REG_ADDR_W-1:0] raddr2 = ifid_valid_cur ? ifid_inst_cur[24:20] : {`REG_ADDR_W{1'b0}};
    wire [`XLEN-1:0] rdata1;
    wire [`XLEN-1:0] rdata2;
    wire wb_we;
    wire [`HART_ID_W-1:0] wb_hart_id;
    wire [`REG_ADDR_W-1:0] waddr;
    wire [`XLEN-1:0] wdata;

    wire [11:0] csr_addr;
    wire csr_we;
    wire [`XLEN-1:0] csr_wdata;
    wire csr_re;
    wire [`XLEN-1:0] csr_rdata;
    wire [`XLEN-1:0] mstatus;
    wire [`XLEN-1:0] mie;
    wire [`XLEN-1:0] mip;
    wire [`XLEN-1:0] mtvec;
    wire [`XLEN-1:0] mepc;
    wire [`XLEN-1:0] mcause;

    wire [`XLEN-1:0] cur_pc = pc[exec_hart];
    wire trap_set_raw;
    wire trap_set;
    wire [`HART_ID_W-1:0] trap_hart_id;
    wire [`XLEN-1:0] trap_vector;
    wire [`XLEN-1:0] trap_mepc;
    wire [`XLEN-1:0] trap_mcause;
    wire trap_mret;

    wire branch_taken;
    wire [`XLEN-1:0] branch_target;
    wire mem_is_data;
    wire ifetch_any_inflight;
    wire mem_req_data;
    wire mem_we_data;
    wire [`ADDR_W-1:0] mem_addr_data;
    wire [`XLEN-1:0] mem_wdata_data;
    wire [`XLEN-1:0] mem_wb_data;
    wire mem_stall;
    wire muldiv_wait;
    wire wb_stall;
    wire pipe_stall;
    wire fetch_block_h0 = exec_valid &&
                          (exec_hart == {`HART_ID_W{1'b0}}) &&
                          (trap_set || trap_mret || branch_taken);
    wire fetch_block_h1 = exec_valid &&
                          (exec_hart == {{(`HART_ID_W-1){1'b0}}, 1'b1}) &&
                          (trap_set || trap_mret || branch_taken);
    wire fetch_pick_h0 = !ifid_valid[0] && !fetch_block_h0;
    wire fetch_pick_h1 = !ifid_valid[1] && !fetch_block_h1 && !fetch_pick_h0;
    wire fetch_any = fetch_pick_h0 || fetch_pick_h1;
    wire fetch_issue = !mem_inflight && fetch_any && !mem_req_data;
    wire [`HART_ID_W-1:0] fetch_hart_sel =
        fetch_pick_h0 ? {`HART_ID_W{1'b0}} : {{(`HART_ID_W-1){1'b0}}, 1'b1};
    wire [`XLEN-1:0] fetch_pc_sel = fetch_pick_h0 ? pc[0] : pc[1];
    wire if_req = ifetch_req || fetch_issue;
    wire [`XLEN-1:0] if_pc_req = ifetch_req ? ifetch_pc_d : fetch_pc_sel;
    wire if_mem_req;
    wire [`ADDR_W-1:0] if_mem_addr;
    wire [`XLEN-1:0] if_inst;
    wire if_inst_valid;
    wire [`XLEN-1:0] if_pc_next;

    wire [`REG_ADDR_W-1:0] id_rs1;
    wire [`REG_ADDR_W-1:0] id_rs2;
    wire [`REG_ADDR_W-1:0] id_rd;
    wire [6:0] id_opcode;
    wire [2:0] id_funct3;
    wire [6:0] id_funct7;
    wire [`XLEN-1:0] id_imm;
    wire [`XLEN-1:0] id_rs1_val;
    wire [`XLEN-1:0] id_rs2_val;

    wire [`XLEN-1:0] ex_alu_result;
    wire ex_branch_taken;
    wire [`XLEN-1:0] ex_branch_target;
    assign branch_taken = idex_valid_cur && ex_branch_taken;
    assign branch_target = ex_branch_target;

    wire ex_is_op_imm = (idex_opcode_cur == 7'b0010011);
    wire ex_is_op     = (idex_opcode_cur == 7'b0110011) && (idex_funct7_cur != 7'b0000001);
    wire ex_is_lui   = (idex_opcode_cur == 7'b0110111);
    wire ex_is_auipc = (idex_opcode_cur == 7'b0010111);
    wire ex_is_jal   = (idex_opcode_cur == 7'b1101111);
    wire ex_is_jalr  = (idex_opcode_cur == 7'b1100111) && (idex_funct3_cur == 3'b000);
    wire ex_is_branch = (idex_opcode_cur == 7'b1100011);
    wire ex_is_load  = (idex_opcode_cur == 7'b0000011) && (idex_funct3_cur == 3'b010);
    wire ex_is_store = (idex_opcode_cur == 7'b0100011) && (idex_funct3_cur == 3'b010);
    wire ex_is_system = (idex_opcode_cur == 7'b1110011);
    wire ex_is_csrrw = ex_is_system && (idex_funct3_cur == 3'b001);
    wire ex_is_csrrs = ex_is_system && (idex_funct3_cur == 3'b010);
    wire ex_is_csr = ex_is_csrrw || ex_is_csrrs;
    wire ex_is_mret = ex_is_system && (idex_funct3_cur == 3'b000) && (idex_inst_cur[31:20] == 12'h302);
    wire ex_is_muldiv = (idex_opcode_cur == 7'b0110011) && (idex_funct7_cur == 7'b0000001);
    reg [2:0] ex_muldiv_op;
    wire ex_mem_op = idex_valid_cur && (ex_is_load || ex_is_store);
    wire ex_wb_en = idex_valid_cur &&
                    (ex_is_op_imm || ex_is_op || ex_is_load || ex_is_csr ||
                     ex_is_lui || ex_is_auipc || ex_is_jal || ex_is_jalr) &&
                    !ex_is_muldiv;
    wire [`REG_ADDR_W-1:0] ex_wb_rd = idex_rd_cur;
    wire [`XLEN-1:0] ex_wb_data_raw = ex_is_csr ? csr_rdata :
                                      (ex_is_jal || ex_is_jalr) ? (idex_pc_cur + 32'd4) :
                                      ex_alu_result;
    wire [`HART_ID_W-1:0] ex_wb_hart_id = idex_hart_id_cur;
    wire muldiv_wb_fire;
    wire [`XLEN-1:0] ex_rs1_val;
    wire [`XLEN-1:0] ex_rs2_val;

    wire muldiv_issue = exec_valid && idex_valid_cur && ex_is_muldiv &&
                        !muldiv_busy && !mem_stall && !wb_stall && !trap_set;
    assign muldiv_wait = exec_valid && idex_valid_cur && ex_is_muldiv && muldiv_busy;

    assign pipe_stall = mem_stall || muldiv_wait || wb_stall;

    always @(*) begin
        ex_muldiv_op = `MULDIV_OP_MUL;
        case (idex_funct3_cur)
            3'b000: ex_muldiv_op = `MULDIV_OP_MUL;
            3'b001: ex_muldiv_op = `MULDIV_OP_MULH;
            3'b010: ex_muldiv_op = `MULDIV_OP_MULHSU;
            3'b011: ex_muldiv_op = `MULDIV_OP_MULHU;
            3'b100: ex_muldiv_op = `MULDIV_OP_DIV;
            3'b101: ex_muldiv_op = `MULDIV_OP_DIVU;
            3'b110: ex_muldiv_op = `MULDIV_OP_REM;
            3'b111: ex_muldiv_op = `MULDIV_OP_REMU;
            default: ex_muldiv_op = `MULDIV_OP_MUL;
        endcase
    end

    always @(*) begin
        blocked_n = blocked;
        if (muldiv_issue) begin
            blocked_n[exec_hart] = 1'b1;
        end
        if (muldiv_wb_fire) begin
            blocked_n[muldiv_pending_hart_id] = 1'b0;
        end
    end

    always @(posedge clk) begin
        if (!rst_n) begin
            blocked <= {`HART_NUM{1'b0}};
        end else begin
            blocked <= blocked_n;
        end
    end

    wire mem_ready_ifetch = cpu_mem_ready && mem_req_d && !mem_is_data_d;
    wire mem_ready_data;

    assign ifetch_any_inflight = ifetch_req;

    always @(posedge clk) begin
        if (!rst_n) begin
            muldiv_pending <= 1'b0;
            muldiv_pending_result <= {`XLEN{1'b0}};
            muldiv_pending_hart_id <= {`HART_ID_W{1'b0}};
            muldiv_pending_rd <= {`REG_ADDR_W{1'b0}};
            ifetch_hart_d <= {`HART_ID_W{1'b0}};
            ifetch_pc_d <= {`XLEN{1'b0}};
            ifetch_req <= 1'b0;
            mem_inflight <= 1'b0;
            mem_inflight_is_data <= 1'b0;
            mem_inflight_addr <= {`ADDR_W{1'b0}};
            mem_inflight_we <= 1'b0;
            mem_inflight_wdata <= {`XLEN{1'b0}};
            mem_req_d <= 1'b0;
            mem_is_data_d <= 1'b0;
            for (h = 0; h < `HART_NUM; h = h + 1) begin
                ifetch_kill[h] <= 1'b0;
            end
        end else begin
            mem_req_d <= mem_inflight;
            mem_is_data_d <= mem_inflight_is_data;
            if (muldiv_done && !muldiv_pending) begin
                muldiv_pending <= 1'b1;
                muldiv_pending_result <= muldiv_result;
                muldiv_pending_hart_id <= muldiv_done_hart_id;
                muldiv_pending_rd <= muldiv_done_rd;
            end else if (muldiv_wb_fire) begin
                muldiv_pending <= 1'b0;
            end

            if (mem_inflight && cpu_mem_ready) begin
                if (!mem_inflight_is_data) begin
                    ifetch_req <= 1'b0;
                    if (ifetch_kill[ifetch_hart_d]) begin
                        ifetch_kill[ifetch_hart_d] <= 1'b0;
                    end
                end
                mem_inflight <= 1'b0;
                mem_inflight_is_data <= 1'b0;
                mem_inflight_we <= 1'b0;
                mem_inflight_wdata <= {`XLEN{1'b0}};
            end

            if (!mem_inflight) begin
                if (mem_req_data) begin
                    mem_inflight <= 1'b1;
                    mem_inflight_is_data <= 1'b1;
                    mem_inflight_addr <= mem_addr_data;
                    mem_inflight_we <= mem_we_data;
                    mem_inflight_wdata <= mem_wdata_data;
                end else if (fetch_issue) begin
                    mem_inflight <= 1'b1;
                    mem_inflight_is_data <= 1'b0;
                    mem_inflight_addr <= fetch_pc_sel;
                    mem_inflight_we <= 1'b0;
                    mem_inflight_wdata <= {`XLEN{1'b0}};
                    ifetch_hart_d <= fetch_hart_sel;
                    ifetch_pc_d <= fetch_pc_sel;
                    ifetch_req <= 1'b1;
                end
            end

            if (exec_valid && !pipe_stall && (trap_set || trap_mret || branch_taken)) begin
                // Drop the next IFetch response for this hart only when a prior fetch is in-flight.
                if (ifetch_req && (ifetch_hart_d == exec_hart) && !mem_ready_ifetch) begin
                    ifetch_kill[exec_hart] <= 1'b1;
                end
            end
        end
    end

    always @(posedge clk) begin
        if (!rst_n) begin
            for (h = 0; h < `HART_NUM; h = h + 1) begin
                pc[h] <= `RESET_VECTOR;
                ifid_valid[h] <= 1'b0;
                ifid_pc[h] <= {`XLEN{1'b0}};
                ifid_inst[h] <= 32'b0;
                idex_valid[h] <= 1'b0;
                idex_pc[h] <= {`XLEN{1'b0}};
                idex_inst[h] <= 32'b0;
                idex_hart_id[h] <= {`HART_ID_W{1'b0}};
                idex_rs1[h] <= {`REG_ADDR_W{1'b0}};
                idex_rs2[h] <= {`REG_ADDR_W{1'b0}};
                idex_rd[h] <= {`REG_ADDR_W{1'b0}};
                idex_opcode[h] <= 7'b0;
                idex_funct3[h] <= 3'b0;
                idex_funct7[h] <= 7'b0;
                idex_imm[h] <= {`XLEN{1'b0}};
                idex_rs1_val[h] <= {`XLEN{1'b0}};
                idex_rs2_val[h] <= {`XLEN{1'b0}};
                exmem_valid[h] <= 1'b0;
                exmem_hart_id[h] <= {`HART_ID_W{1'b0}};
                exmem_rd[h] <= {`REG_ADDR_W{1'b0}};
                exmem_alu_result[h] <= {`XLEN{1'b0}};
                exmem_rs2_val[h] <= {`XLEN{1'b0}};
                exmem_is_load[h] <= 1'b0;
                exmem_mem_we[h] <= 1'b0;
                exmem_wb_en[h] <= 1'b0;
                exmem_wb_data_raw[h] <= {`XLEN{1'b0}};
                exwb_valid[h] <= 1'b0;
                exwb_hart_id[h] <= {`HART_ID_W{1'b0}};
                exwb_rd[h] <= {`REG_ADDR_W{1'b0}};
                exwb_data[h] <= {`XLEN{1'b0}};
            end
        end else begin
            if (ifetch_req && mem_ready_ifetch) begin
                if (!ifetch_kill[ifetch_hart_d] &&
                    !(ifetch_hart_d == exec_hart &&
                      (trap_set || trap_mret || branch_taken))) begin
                    ifid_valid[ifetch_hart_d] <= 1'b1;
                    ifid_pc[ifetch_hart_d] <= ifetch_pc_d;
                    ifid_inst[ifetch_hart_d] <= if_inst;
                    pc[ifetch_hart_d] <= ifetch_pc_d + 32'd4;
                end
            end

            if (exec_valid) begin
                if (!pipe_stall) begin
                    if (trap_set) begin
                    exmem_valid[exec_hart] <= 1'b0;
                    exmem_is_load[exec_hart] <= 1'b0;
                    exmem_mem_we[exec_hart] <= 1'b0;
                    exmem_wb_en[exec_hart] <= 1'b0;
                    exwb_valid[exec_hart] <= 1'b0;
                end else begin
                    exwb_valid[exec_hart] <= exmem_wb_en_cur;
                    exwb_hart_id[exec_hart] <= exmem_hart_id_cur;
                    exwb_rd[exec_hart] <= exmem_rd_cur;
                    exwb_data[exec_hart] <= mem_wb_data;

                    exmem_valid[exec_hart] <= idex_valid_cur && (ex_wb_en || ex_mem_op);
                    exmem_hart_id[exec_hart] <= ex_wb_hart_id;
                    exmem_rd[exec_hart] <= ex_wb_rd;
                    exmem_alu_result[exec_hart] <= ex_alu_result;
                    exmem_rs2_val[exec_hart] <= ex_rs2_val;
                    exmem_is_load[exec_hart] <= ex_is_load;
                    exmem_mem_we[exec_hart] <= ex_is_store;
                    exmem_wb_en[exec_hart] <= ex_wb_en;
                    exmem_wb_data_raw[exec_hart] <= ex_wb_data_raw;
                end
                end

                if (trap_set) begin
                    pc[exec_hart] <= trap_vector;
                    ifid_valid[exec_hart] <= 1'b0;
                    idex_valid[exec_hart] <= 1'b0;
                end else if (trap_mret) begin
                    pc[exec_hart] <= mepc;
                    ifid_valid[exec_hart] <= 1'b0;
                    idex_valid[exec_hart] <= 1'b0;
                end else if (branch_taken) begin
                    pc[exec_hart] <= branch_target;
                    ifid_valid[exec_hart] <= 1'b0;
                    idex_valid[exec_hart] <= 1'b0;
                end else begin
                    if (ifid_valid[exec_hart]) begin
                        idex_valid[exec_hart] <= 1'b1;
                        idex_pc[exec_hart] <= ifid_pc[exec_hart];
                        idex_inst[exec_hart] <= ifid_inst[exec_hart];
                        idex_hart_id[exec_hart] <= exec_hart;
                        idex_rs1[exec_hart] <= id_rs1;
                        idex_rs2[exec_hart] <= id_rs2;
                        idex_rd[exec_hart] <= id_rd;
                        idex_opcode[exec_hart] <= id_opcode;
                        idex_funct3[exec_hart] <= id_funct3;
                        idex_funct7[exec_hart] <= id_funct7;
                        idex_imm[exec_hart] <= id_imm;
                        idex_rs1_val[exec_hart] <= id_rs1_val;
                        idex_rs2_val[exec_hart] <= id_rs2_val;
                    end else begin
                        idex_valid[exec_hart] <= 1'b0;
                    end
                end

                if (!pipe_stall && !trap_set && !trap_mret && !branch_taken) begin
                    if (ifid_valid[exec_hart] &&
                        !(ifetch_req && mem_ready_ifetch &&
                          (ifetch_hart_d == exec_hart))) begin
                        ifid_valid[exec_hart] <= 1'b0;
                    end
                end
            end
        end
    end

    barrel_sched u_sched (
        .clk(clk),
        .rst_n(rst_n),
        .blocked(blocked),
        .hold(mem_stall),
        .cur_hart(cur_hart),
        .cur_valid(cur_valid)
    );

    regfile_bank u_regfile (
        .clk(clk),
        .rst_n(rst_n),
        .r_hart_id(exec_hart),
        .raddr1(raddr1),
        .raddr2(raddr2),
        .rdata1(rdata1),
        .rdata2(rdata2),
        .w_en(wb_we),
        .w_hart_id(wb_hart_id),
        .waddr(waddr),
        .wdata(wdata)
    );

    csr_file u_csr (
        .clk(clk),
        .rst_n(rst_n),
        .hart_id(exec_hart),
        .csr_addr(csr_addr),
        .csr_we(csr_we),
        .csr_wdata(csr_wdata),
        .csr_re(csr_re),
        .csr_rdata(csr_rdata),
        .ext_irq(ext_irq),
        .trap_set(trap_set),
        .trap_hart_id(trap_hart_id),
        .trap_mepc(trap_mepc),
        .trap_mcause(trap_mcause),
        .trap_mret(trap_mret),
        .mstatus_o(mstatus),
        .mie_o(mie),
        .mip_o(mip),
        .mtvec_o(mtvec),
        .mepc_o(mepc),
        .mcause_o(mcause)
    );

    trap_ctrl u_trap (
        .clk(clk),
        .rst_n(rst_n),
        .hart_id(exec_hart),
        .pc_in(cur_pc),
        .mtvec(mtvec),
        .mstatus(mstatus),
        .mie(mie),
        .mip(mip),
        .take_trap(trap_set_raw),
        .trap_hart_id(trap_hart_id),
        .trap_vector(trap_vector),
        .trap_mepc(trap_mepc),
        .trap_mcause(trap_mcause)
    );

    if_stage u_if (
        .pc_in(if_pc_req),
        .if_valid(if_req),
        .mem_rdata(cpu_mem_rdata),
        .mem_ready(cpu_mem_ready),
        .mem_req(if_mem_req),
        .mem_addr(if_mem_addr),
        .inst_out(if_inst),
        .inst_valid(if_inst_valid),
        .pc_next(if_pc_next)
    );

    id_stage u_id (
        .inst_in(ifid_inst_cur),
        .pc_in(ifid_pc_cur),
        .rdata1(rdata1),
        .rdata2(rdata2),
        .rs1(id_rs1),
        .rs2(id_rs2),
        .rd(id_rd),
        .opcode(id_opcode),
        .funct3(id_funct3),
        .funct7(id_funct7),
        .imm(id_imm),
        .rs1_val(id_rs1_val),
        .rs2_val(id_rs2_val)
    );

    hazard_fwd u_fwd (
        .rs1_addr(idex_rs1_cur),
        .rs2_addr(idex_rs2_cur),
        .rs1_val_in(idex_rs1_val_cur),
        .rs2_val_in(idex_rs2_val_cur),
        .exmem_wb_en(exmem_wb_en_cur),
        .exmem_rd(exmem_rd_cur),
        .exmem_wb_data(mem_wb_data),
        .exwb_wb_en(exwb_valid_cur),
        .exwb_rd(exwb_rd_cur),
        .exwb_wb_data(exwb_data_cur),
        .rs1_val_out(ex_rs1_val),
        .rs2_val_out(ex_rs2_val)
    );

    assign mem_ready_data = cpu_mem_ready && mem_req_d && mem_is_data_d;

    mem_stage u_mem (
        .exmem_valid(exmem_valid_cur && exec_valid),
        .exmem_is_load(exmem_is_load_cur),
        .exmem_mem_we(exmem_mem_we_cur),
        .exmem_addr(exmem_alu_result_cur),
        .exmem_wdata(exmem_rs2_val_cur),
        .exmem_wb_data_raw(exmem_wb_data_raw_cur),
        .mem_ready(mem_ready_data),
        .mem_rdata(cpu_mem_rdata),
        .mem_req(mem_req_data),
        .mem_we(mem_we_data),
        .mem_addr(mem_addr_data),
        .mem_wdata(mem_wdata_data),
        .mem_wb_data(mem_wb_data),
        .mem_stall(mem_stall)
    );

    wb_stage u_wb (
        .exec_valid(exec_valid),
        .mem_stall(mem_stall),
        .exwb_valid(exwb_valid_cur),
        .exwb_hart_id(exwb_hart_id_cur),
        .exwb_rd(exwb_rd_cur),
        .exwb_data(exwb_data_cur),
        .muldiv_pending(muldiv_pending),
        .muldiv_pending_hart_id(muldiv_pending_hart_id),
        .muldiv_pending_rd(muldiv_pending_rd),
        .muldiv_pending_result(muldiv_pending_result),
        .wb_we(wb_we),
        .wb_hart_id(wb_hart_id),
        .wb_rd(waddr),
        .wb_data(wdata),
        .wb_stall(wb_stall),
        .muldiv_wb_fire(muldiv_wb_fire)
    );

    ex_stage u_ex (
        .opcode(idex_opcode_cur),
        .funct3(idex_funct3_cur),
        .funct7(idex_funct7_cur),
        .rs1_val(ex_rs1_val),
        .rs2_val(ex_rs2_val),
        .imm(idex_imm_cur),
        .pc_in(idex_pc_cur),
        .alu_result(ex_alu_result),
        .branch_taken(ex_branch_taken),
        .branch_target(ex_branch_target)
    );

    assign trap_set = trap_set_raw && exec_valid && !pipe_stall;
    assign trap_mret = ex_is_mret && exec_valid && !pipe_stall;

    assign csr_addr = idex_inst_cur[31:20];
    assign csr_re = ex_is_csr && exec_valid && !pipe_stall;
    assign csr_wdata = ex_is_csrrw ? ex_rs1_val : (csr_rdata | ex_rs1_val);
    assign csr_we = ex_is_csr && exec_valid && !pipe_stall &&
                    (ex_is_csrrw || (ex_is_csrrs && (idex_rs1_cur != {`REG_ADDR_W{1'b0}})));

    assign mem_is_data = mem_inflight && mem_inflight_is_data;
    assign cpu_mem_req   = mem_inflight;
    assign cpu_mem_we    = mem_inflight && mem_inflight_is_data && mem_inflight_we;
    assign cpu_mem_addr  = mem_inflight ? mem_inflight_addr : {`ADDR_W{1'b0}};
    assign cpu_mem_wdata = mem_inflight ? mem_inflight_wdata : {`XLEN{1'b0}};

    assign muldiv_start   = muldiv_issue;
    assign muldiv_op      = ex_muldiv_op;
    assign muldiv_a       = ex_rs1_val;
    assign muldiv_b       = ex_rs2_val;
    assign muldiv_hart_id = idex_hart_id_cur;
    assign muldiv_rd      = idex_rd_cur;
endmodule
