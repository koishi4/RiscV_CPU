`include "defines.vh"

module wb_stage(
    input clk,
    input rst_n
);
    // TODO: writeback stage.
endmodule
