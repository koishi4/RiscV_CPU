`include "defines.vh"

module id_stage(
    input clk,
    input rst_n
);
    // TODO: decode/register fetch stage.
endmodule
