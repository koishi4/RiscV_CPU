`include "defines.vh"

module csr_file(
    input clk,
    input rst_n
);
    // TODO: per-hart CSR storage and access.
endmodule
