`include "defines.vh"

module mem_stage(
    input clk,
    input rst_n
);
    // TODO: memory access stage.
endmodule
