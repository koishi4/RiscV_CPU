`include "defines.vh"

module if_stage(
    input clk,
    input rst_n
);
    // TODO: instruction fetch stage.
endmodule
