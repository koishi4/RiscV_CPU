`include "defines.vh"

module hazard_fwd(
    input clk,
    input rst_n
);
    // TODO: hazard detection and forwarding.
endmodule
